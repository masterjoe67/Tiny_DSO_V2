PLL_Master_inst : PLL_Master PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig,
		c1	 => c1_sig
	);
